module (
    clk,
    rst,
    addr,
    VRAM_available,
    color_in
);











endmodule