module control_paint(
    clk,
    rst,
    in_init,
    w_C,
    w_Enter,
    x_out,
    y_out,
    in_C,
    paleta,
    pixel_data,
    paint,
    selector,
    out_PAINT,
    out_DRAW_CURSOR,
    out_CURSOR_PALETA,

);

endmodule