module BCD(
    clk,
    rst,
    init,
    in_BIN,
    out_UND,
    out_DEC,
    out_CEN,
    out_DONE  
);
input rst;
input clk;
input init;
input in_BIN;

    
endmodule //BCD

